module controller (
	iClk,
	iPSR,
	iInstruction,
	opc,
	oALU_source1,
	oALU_source2
);


endmodule